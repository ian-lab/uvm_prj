`ifndef MY_MODEL_SV
`define MY_MODEL_SV

import uvm_pkg::*;
`include "uvm_macros.svh"
`include "my_transaction.sv"

class my_model extends uvm_component;
    `uvm_component_utils(my_model)

    uvm_blocking_get_port #(my_trans) port;
    uvm_analysis_port #(my_trans) ap;

    function new(string name="my_model", uvm_component parent);
        super.new(name, parent);
    endfunction 

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        port = new("port",this);
        ap = new("ap",this);
    endfunction

    task main_phase(uvm_phase phase);
        my_trans tr;
        my_trans new_tr;
        int message_frame, t;
        bit [31:0] w_seq [$];
        bit [63:0] message_seq [$];
        bit [31:0] H0,H1,H2,H3,H4,A,B,C,D,E,temp,k,f,w;
        bit [63:0] andmask, ormask, pad_one;
        bit [ 2:0] zero_pad_len; 
        bit [63:0] len_pad;
        bit [63:0] pad_message_len;
        bit [159:0] hash;
        while(1) begin
            port.get(tr);
            new_tr = new("new_tr");
            new_tr.copy(tr);
            message_seq.delete();

            //data
            foreach(tr.drv_data[i]) begin
                message_seq.push_back(tr.drv_data[i]);
            end
            // pad one
            if(tr.drv_len % 64==0) begin
                pad_one = {1'b1, {63{1'b0}}};
                message_seq.push_back(pad_one );
            end
            else begin
                pad_one = message_seq.pop_back();
                andmask = Andmask(tr.drv_len);
                ormask = Ormask(tr.drv_len);
                pad_one = (pad_one & andmask) | ormask;
                message_seq.push_back(pad_one);
            end
            // pad zero
            zero_pad_len = 8 - tr.drv_len[63:6] % 8 - 1 - 1 ;
            for(int a = 0; a < zero_pad_len; a=a+1)
                message_seq.push_back(64'b0);
            // pad len
            len_pad = 64'b0 | tr.drv_len;
            message_seq.push_back(len_pad);
            pad_message_len = tr.drv_len + (512-(tr.drv_len+64)%512) + 64;
            H0 = 32'h67452301; H1 = 32'hEFCDAB89;
            H2 = 32'h98BADCFE; H3 = 32'h10325476;
            H4 = 32'hC3D2E1F0;
            // foreach(message_seq[i]) begin
            //     `uvm_info(get_type_name(), $sformatf("data is 'h%16x", message_seq[i]), UVM_LOW)
            // end
            for (message_frame=0; message_frame<(pad_message_len/512); message_frame=message_frame+1)begin
                A = H0; B = H1; C = H2; D = H3; E = H4;
                for (t=0; t<80; t=t+1)begin
                    if(t < 16) begin
                        w_seq[0]  = message_seq[message_frame*8][63:32];
                        w_seq[1]  = message_seq[message_frame*8][31:0];
                        w_seq[2]  = message_seq[message_frame*8+1][63:32];
                        w_seq[3]  = message_seq[message_frame*8+1][31:0];
                        w_seq[4]  = message_seq[message_frame*8+2][63:32];
                        w_seq[5]  = message_seq[message_frame*8+2][31:0];
                        w_seq[6]  = message_seq[message_frame*8+3][63:32];
                        w_seq[7]  = message_seq[message_frame*8+3][31:0];
                        w_seq[8]  = message_seq[message_frame*8+4][63:32];
                        w_seq[9]  = message_seq[message_frame*8+4][31:0];
                        w_seq[10] = message_seq[message_frame*8+5][63:32];
                        w_seq[11] = message_seq[message_frame*8+5][31:0];
                        w_seq[12] = message_seq[message_frame*8+6][63:32];
                        w_seq[13] = message_seq[message_frame*8+6][31:0];
                        w_seq[14] = message_seq[message_frame*8+7][63:32];
                        w_seq[15] = message_seq[message_frame*8+7][31:0];
                        w = w_seq[t];
                    end
                    else begin
                        w = w_seq[13] ^ w_seq[8] ^ w_seq[2] ^ w_seq[0];
                        w = {w[30:0], w[31]};
                        w_seq.push_back(w);
                       void'(w_seq.pop_front());
                    end
                       
                    if (t <= 19)begin
                        k = 64'h5A827999;
                        f = (B & C) | (~B & D);
                    end
                    else if (t>=20 && t<=39)begin
                        k = 64'h6ED9EBA1;
                        f = B ^ C ^ D;
                    end
                    else if (t>=40 && t<=59)begin
                        k = 64'h8F1BBCDC;
                        f = (B & C) | (B & D) | (C & D);
                    end
                    else if (t>=60 && t<=79)begin
                        k = 64'hCA62C1D6;
                        f = B ^ C ^ D;
                    end
                    temp ={A[26:0], A[31:27]} + f + E + w + k;
                   
                    E = D;
                    D = C;
                    C = {B[1:0], B[31:2]};
                    B = A;
                    A = temp;
                    // `uvm_info(get_type_name(), $sformatf("t is 'h%2d",t+1), UVM_LOW)
                    // `uvm_info(get_type_name(), $sformatf("w is 'h%8x",w), UVM_LOW)
                    //  `uvm_info(get_type_name(), $sformatf("A is 'h%8x",A), UVM_LOW)
                    // `uvm_info(get_type_name(), $sformatf("B is 'h%8x",B), UVM_LOW)
                    // `uvm_info(get_type_name(), $sformatf("c is 'h%8x",C), UVM_LOW)
                    // `uvm_info(get_type_name(), $sformatf("d is 'h%8x",D), UVM_LOW)
                    // `uvm_info(get_type_name(), $sformatf("e is 'h%8x",E), UVM_LOW)
                    // `uvm_info(get_type_name(), $sformatf("F is 'h%8x",f), UVM_LOW)
                    // `uvm_info(get_type_name(), $sformatf("k is 'h%8x",k), UVM_LOW)
                    if (t == 7'd79) begin
                        H0 = H0 + A;
                        H1 = H1 + B;
                        H2 = H2 + C;
                        H3 = H3 + D;
                        H4 = H4 + E;
                    end
                    hash = {H0, H1, H2, H3, H4};
                end
            end
            new_tr.hash = hash;
            // `uvm_info(get_type_name(), $sformatf("hash is 'h%40x", hash), UVM_LOW)
            ap.write(new_tr);
        end
    endtask 

    function bit[63:0] Andmask(bit[64:0] data);
        case(data[5:0])
            6'd0:   return 64'b1000000000000000000000000000000000000000000000000000000000000000;
		    6'd1:   return 64'b1100000000000000000000000000000000000000000000000000000000000000;
		    6'd2:   return 64'b1110000000000000000000000000000000000000000000000000000000000000;
		    6'd3:   return 64'b1111000000000000000000000000000000000000000000000000000000000000;
		    6'd4:   return 64'b1111100000000000000000000000000000000000000000000000000000000000;
		    6'd5:   return 64'b1111110000000000000000000000000000000000000000000000000000000000;
		    6'd6:   return 64'b1111111000000000000000000000000000000000000000000000000000000000;
		    6'd7:   return 64'b1111111100000000000000000000000000000000000000000000000000000000;
		    6'd8:   return 64'b1111111110000000000000000000000000000000000000000000000000000000;
		    6'd9:   return 64'b1111111111000000000000000000000000000000000000000000000000000000;
		    6'd10:  return 64'b1111111111100000000000000000000000000000000000000000000000000000;
		    6'd11:  return 64'b1111111111110000000000000000000000000000000000000000000000000000;
		    6'd12:  return 64'b1111111111111000000000000000000000000000000000000000000000000000;
		    6'd13:  return 64'b1111111111111100000000000000000000000000000000000000000000000000;
		    6'd14:  return 64'b1111111111111110000000000000000000000000000000000000000000000000;
		    6'd15:  return 64'b1111111111111111000000000000000000000000000000000000000000000000;
		    6'd16:  return 64'b1111111111111111100000000000000000000000000000000000000000000000;
		    6'd17:  return 64'b1111111111111111110000000000000000000000000000000000000000000000;
		    6'd18:  return 64'b1111111111111111111000000000000000000000000000000000000000000000;
		    6'd19:  return 64'b1111111111111111111100000000000000000000000000000000000000000000;
		    6'd20:  return 64'b1111111111111111111110000000000000000000000000000000000000000000;
		    6'd21:  return 64'b1111111111111111111111000000000000000000000000000000000000000000;
		    6'd22:  return 64'b1111111111111111111111100000000000000000000000000000000000000000;
		    6'd23:  return 64'b1111111111111111111111110000000000000000000000000000000000000000;
		    6'd24:  return 64'b1111111111111111111111111000000000000000000000000000000000000000;
		    6'd25:  return 64'b1111111111111111111111111100000000000000000000000000000000000000;
		    6'd26:  return 64'b1111111111111111111111111110000000000000000000000000000000000000;
		    6'd27:  return 64'b1111111111111111111111111111000000000000000000000000000000000000;
		    6'd28:  return 64'b1111111111111111111111111111100000000000000000000000000000000000;
		    6'd29:  return 64'b1111111111111111111111111111110000000000000000000000000000000000;
		    6'd30:  return 64'b1111111111111111111111111111111000000000000000000000000000000000;
		    6'd31:  return 64'b1111111111111111111111111111111100000000000000000000000000000000;
		    6'd32:  return 64'b1111111111111111111111111111111110000000000000000000000000000000;
		    6'd33:  return 64'b1111111111111111111111111111111111000000000000000000000000000000;
		    6'd34:  return 64'b1111111111111111111111111111111111100000000000000000000000000000;
		    6'd35:  return 64'b1111111111111111111111111111111111110000000000000000000000000000;
		    6'd36:  return 64'b1111111111111111111111111111111111111000000000000000000000000000;
		    6'd37:  return 64'b1111111111111111111111111111111111111100000000000000000000000000;
		    6'd38:  return 64'b1111111111111111111111111111111111111110000000000000000000000000;
		    6'd39:  return 64'b1111111111111111111111111111111111111111000000000000000000000000;
		    6'd40:  return 64'b1111111111111111111111111111111111111111100000000000000000000000;
		    6'd41:  return 64'b1111111111111111111111111111111111111111110000000000000000000000;
		    6'd42:  return 64'b1111111111111111111111111111111111111111111000000000000000000000;
		    6'd43:  return 64'b1111111111111111111111111111111111111111111100000000000000000000;
		    6'd44:  return 64'b1111111111111111111111111111111111111111111110000000000000000000;
		    6'd45:  return 64'b1111111111111111111111111111111111111111111111000000000000000000;
		    6'd46:  return 64'b1111111111111111111111111111111111111111111111100000000000000000;
		    6'd47:  return 64'b1111111111111111111111111111111111111111111111110000000000000000;
		    6'd48:  return 64'b1111111111111111111111111111111111111111111111111000000000000000;
		    6'd49:  return 64'b1111111111111111111111111111111111111111111111111100000000000000;
		    6'd50:  return 64'b1111111111111111111111111111111111111111111111111110000000000000;
		    6'd51:  return 64'b1111111111111111111111111111111111111111111111111111000000000000;
		    6'd52:  return 64'b1111111111111111111111111111111111111111111111111111100000000000;
		    6'd53:  return 64'b1111111111111111111111111111111111111111111111111111110000000000;
		    6'd54:  return 64'b1111111111111111111111111111111111111111111111111111111000000000;
		    6'd55:  return 64'b1111111111111111111111111111111111111111111111111111111100000000;
		    6'd56:  return 64'b1111111111111111111111111111111111111111111111111111111110000000;
		    6'd57:  return 64'b1111111111111111111111111111111111111111111111111111111111000000;
		    6'd58:  return 64'b1111111111111111111111111111111111111111111111111111111111100000;
		    6'd59:  return 64'b1111111111111111111111111111111111111111111111111111111111110000;
		    6'd60:  return 64'b1111111111111111111111111111111111111111111111111111111111111000;
		    6'd61:  return 64'b1111111111111111111111111111111111111111111111111111111111111100;
		    6'd62:  return 64'b1111111111111111111111111111111111111111111111111111111111111110;
		    6'd63:  return 64'b1111111111111111111111111111111111111111111111111111111111111111;
	    endcase
    endfunction

    function bit[63:0] Ormask(bit[64:0] data);
        case(data[5:0])
            6'd0:   return 64'b1000000000000000000000000000000000000000000000000000000000000000;
		    6'd1:   return 64'b0100000000000000000000000000000000000000000000000000000000000000;
		    6'd2:   return 64'b0010000000000000000000000000000000000000000000000000000000000000;
		    6'd3:   return 64'b0001000000000000000000000000000000000000000000000000000000000000;
		    6'd4:   return 64'b0000100000000000000000000000000000000000000000000000000000000000;
		    6'd5:   return 64'b0000010000000000000000000000000000000000000000000000000000000000;
		    6'd6:   return 64'b0000001000000000000000000000000000000000000000000000000000000000;
		    6'd7:   return 64'b0000000100000000000000000000000000000000000000000000000000000000;
		    6'd8:   return 64'b0000000010000000000000000000000000000000000000000000000000000000;
		    6'd9:   return 64'b0000000001000000000000000000000000000000000000000000000000000000;
		    6'd10:  return 64'b0000000000100000000000000000000000000000000000000000000000000000;
		    6'd11:  return 64'b0000000000010000000000000000000000000000000000000000000000000000;
		    6'd12:  return 64'b0000000000001000000000000000000000000000000000000000000000000000;
		    6'd13:  return 64'b0000000000000100000000000000000000000000000000000000000000000000;
		    6'd14:  return 64'b0000000000000010000000000000000000000000000000000000000000000000;
		    6'd15:  return 64'b0000000000000001000000000000000000000000000000000000000000000000;
		    6'd16:  return 64'b0000000000000000100000000000000000000000000000000000000000000000;
		    6'd17:  return 64'b0000000000000000010000000000000000000000000000000000000000000000;
		    6'd18:  return 64'b0000000000000000001000000000000000000000000000000000000000000000;
		    6'd19:  return 64'b0000000000000000000100000000000000000000000000000000000000000000;
		    6'd20:  return 64'b0000000000000000000010000000000000000000000000000000000000000000;
		    6'd21:  return 64'b0000000000000000000001000000000000000000000000000000000000000000;
		    6'd22:  return 64'b0000000000000000000000100000000000000000000000000000000000000000;
		    6'd23:  return 64'b0000000000000000000000010000000000000000000000000000000000000000;
		    6'd24:  return 64'b0000000000000000000000001000000000000000000000000000000000000000;
		    6'd25:  return 64'b0000000000000000000000000100000000000000000000000000000000000000;
		    6'd26:  return 64'b0000000000000000000000000010000000000000000000000000000000000000;
		    6'd27:  return 64'b0000000000000000000000000001000000000000000000000000000000000000;
		    6'd28:  return 64'b0000000000000000000000000000100000000000000000000000000000000000;
		    6'd29:  return 64'b0000000000000000000000000000010000000000000000000000000000000000;
		    6'd30:  return 64'b0000000000000000000000000000001000000000000000000000000000000000;
		    6'd31:  return 64'b0000000000000000000000000000000100000000000000000000000000000000;
		    6'd32:  return 64'b0000000000000000000000000000000010000000000000000000000000000000;
		    6'd33:  return 64'b0000000000000000000000000000000001000000000000000000000000000000;
		    6'd34:  return 64'b0000000000000000000000000000000000100000000000000000000000000000;
		    6'd35:  return 64'b0000000000000000000000000000000000010000000000000000000000000000;
		    6'd36:  return 64'b0000000000000000000000000000000000001000000000000000000000000000;
		    6'd37:  return 64'b0000000000000000000000000000000000000100000000000000000000000000;
		    6'd38:  return 64'b0000000000000000000000000000000000000010000000000000000000000000;
		    6'd39:  return 64'b0000000000000000000000000000000000000001000000000000000000000000;
		    6'd40:  return 64'b0000000000000000000000000000000000000000100000000000000000000000;
		    6'd41:  return 64'b0000000000000000000000000000000000000000010000000000000000000000;
		    6'd42:  return 64'b0000000000000000000000000000000000000000001000000000000000000000;
		    6'd43:  return 64'b0000000000000000000000000000000000000000000100000000000000000000;
		    6'd44:  return 64'b0000000000000000000000000000000000000000000010000000000000000000;
		    6'd45:  return 64'b0000000000000000000000000000000000000000000001000000000000000000;
		    6'd46:  return 64'b0000000000000000000000000000000000000000000000100000000000000000;
		    6'd47:  return 64'b0000000000000000000000000000000000000000000000010000000000000000;
		    6'd48:  return 64'b0000000000000000000000000000000000000000000000001000000000000000;
		    6'd49:  return 64'b0000000000000000000000000000000000000000000000000100000000000000;
		    6'd50:  return 64'b0000000000000000000000000000000000000000000000000010000000000000;
		    6'd51:  return 64'b0000000000000000000000000000000000000000000000000001000000000000;
		    6'd52:  return 64'b0000000000000000000000000000000000000000000000000000100000000000;
		    6'd53:  return 64'b0000000000000000000000000000000000000000000000000000010000000000;
		    6'd54:  return 64'b0000000000000000000000000000000000000000000000000000001000000000;
		    6'd55:  return 64'b0000000000000000000000000000000000000000000000000000000100000000;
		    6'd56:  return 64'b0000000000000000000000000000000000000000000000000000000010000000;
		    6'd57:  return 64'b0000000000000000000000000000000000000000000000000000000001000000;
		    6'd58:  return 64'b0000000000000000000000000000000000000000000000000000000000100000;
		    6'd59:  return 64'b0000000000000000000000000000000000000000000000000000000000010000;
		    6'd60:  return 64'b0000000000000000000000000000000000000000000000000000000000001000;
		    6'd61:  return 64'b0000000000000000000000000000000000000000000000000000000000000100;
		    6'd62:  return 64'b0000000000000000000000000000000000000000000000000000000000000010;
		    6'd63:  return 64'b0000000000000000000000000000000000000000000000000000000000000001;
	    endcase
    endfunction
endclass 


`endif 