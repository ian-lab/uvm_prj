//=======================================
// module name: sha-1
// author: fan yingbao
// input
//      clk
//      rst_n
//      data_in 
//      valid_in 
//        out_ready   
// output
//      data_pad
//      valid_out
//      in_ready
//=======================================

module message_padder (
    input        clk,
    input        rst_n,
    input [63:0] data_in,
    input        valid_in,
    input        out_ready,

    output reg        valid_out,
    output reg [63:0] data_pad,
    output reg last_block
    
);
localparam LOADLENGTH   = 2'b00;
localparam LOADWORDS    = 2'b01;
localparam PAD_ZERO     = 2'b10;
localparam PAD_LENGTH   = 2'b11;
reg [1:0] state, next_state;

reg  [63:0] message_length;       // length of message       1 bit
reg  [57:0] words_left;           // remaining words        64 bit
reg  [ 2:0] zero_pad_length;      // number of zero-padded  64 bit
reg  [63:0] andMask;
reg  [63:0] orMask;
wire [63:0] data_mask = (data_in & andMask) | orMask; // one-pad

always @(posedge clk or negedge rst_n) begin
    if(!rst_n)begin
        state <= LOADLENGTH;
    end
    else begin
        state <= next_state;
    end
end

always @(posedge clk or negedge rst_n) begin
    if(!rst_n)begin
        message_length <= 64'b0;
        words_left <= 58'b0;
        zero_pad_length = 4'b0;
        data_pad <= 64'b0;
        valid_out <= 1'b0;
        last_block <= 1'b0;
    end
    else begin
        case(state)
            LOADLENGTH : begin
                valid_out <= 1'b0;
                last_block <= 1'b0;
                data_pad <= 64'b0;
                message_length <= data_in;
                words_left <= data_in[63:6];                         // word_left = data_in / 64
                zero_pad_length <= 8 - data_in[63:6] % 8 - 1 - 1 ;   // zero pad = 8 - (message_length/64)%8 - pad one - pad length
            end
            LOADWORDS : begin
                last_block <= 1'b0;
                // if(out_ready && (((message_length[5:0] != 6'd0 | words_left != 58'd0) && valid_in) | (message_length[5:0] == 6'd0 && words_left == 58'd0)))begin
                if(out_ready && ( valid_in | (message_length[5:0] == 6'd0 && words_left == 58'd0)))begin
                    valid_out <= 1'b1;
                    if(words_left == 58'b0)begin
                        data_pad <= data_mask;
                        words_left <= words_left;
                    end
                    else begin
                        data_pad <= data_in;
                        words_left <= words_left - 1'b1;
                    end
                end    
                else begin
                    valid_out <= 1'b0;
                    data_pad <= 64'd0;
                    words_left <= words_left;
                end
            end
            PAD_ZERO :begin
                last_block <= 1'b0;
                if(out_ready) begin
                    valid_out <= 1'b1;
                    zero_pad_length <= zero_pad_length - 1'b1; 
                end
                else
                    valid_out <= 1'b0;
                data_pad = 64'b0;
            end
            PAD_LENGTH : begin
                valid_out <= 1'b1;
                last_block <= 1'b1;
                data_pad <= message_length;
            end
            default: begin
                message_length <= 64'b0;
                words_left <= 58'b0;
                    zero_pad_length = 4'b0;
                data_pad <= 64'b0;
                valid_out <= 1'b0;
                last_block <= 1'b0;
            end
        endcase
    end
end

always @(*) begin
    if(!rst_n)begin
        next_state  = LOADLENGTH;
    end
    else begin
        case(state)
            LOADLENGTH: begin
                if(valid_in)begin
                    next_state = LOADWORDS;
                end
                else begin
                    next_state = LOADLENGTH;
                end
            end
            LOADWORDS: begin
                if(words_left == 58'd0 && out_ready && (valid_in | message_length[5:0] == 0))begin
                    if(zero_pad_length == 64'b0) begin
                        next_state = PAD_LENGTH;
                    end
                    else begin
                        next_state = PAD_ZERO;
                    end
                end
                else begin
                    next_state = LOADWORDS ;
                end
            end
            PAD_ZERO: begin
                if (zero_pad_length == 64'b1)begin
                    next_state = PAD_LENGTH;
                end
                else begin
                    next_state = PAD_ZERO;
                end
            end
            PAD_LENGTH : begin
                next_state = LOADLENGTH;
            end
            default : begin
                next_state = LOADLENGTH;
            end
        endcase
    end
end

always @(*) begin
    case( message_length[5:0] )
        6'd0:   andMask = 64'b1000000000000000000000000000000000000000000000000000000000000000;
        6'd1:   andMask = 64'b1100000000000000000000000000000000000000000000000000000000000000;
        6'd2:   andMask = 64'b1110000000000000000000000000000000000000000000000000000000000000;
        6'd3:   andMask = 64'b1111000000000000000000000000000000000000000000000000000000000000;
        6'd4:   andMask = 64'b1111100000000000000000000000000000000000000000000000000000000000;
        6'd5:   andMask = 64'b1111110000000000000000000000000000000000000000000000000000000000;
        6'd6:   andMask = 64'b1111111000000000000000000000000000000000000000000000000000000000;
        6'd7:   andMask = 64'b1111111100000000000000000000000000000000000000000000000000000000;
        6'd8:   andMask = 64'b1111111110000000000000000000000000000000000000000000000000000000;
        6'd9:   andMask = 64'b1111111111000000000000000000000000000000000000000000000000000000;
        6'd10:  andMask = 64'b1111111111100000000000000000000000000000000000000000000000000000;
        6'd11:  andMask = 64'b1111111111110000000000000000000000000000000000000000000000000000;
        6'd12:  andMask = 64'b1111111111111000000000000000000000000000000000000000000000000000;
        6'd13:  andMask = 64'b1111111111111100000000000000000000000000000000000000000000000000;
        6'd14:  andMask = 64'b1111111111111110000000000000000000000000000000000000000000000000;
        6'd15:  andMask = 64'b1111111111111111000000000000000000000000000000000000000000000000;
        6'd16:  andMask = 64'b1111111111111111100000000000000000000000000000000000000000000000;
        6'd17:  andMask = 64'b1111111111111111110000000000000000000000000000000000000000000000;
        6'd18:  andMask = 64'b1111111111111111111000000000000000000000000000000000000000000000;
        6'd19:  andMask = 64'b1111111111111111111100000000000000000000000000000000000000000000;
        6'd20:  andMask = 64'b1111111111111111111110000000000000000000000000000000000000000000;
        6'd21:  andMask = 64'b1111111111111111111111000000000000000000000000000000000000000000;
        6'd22:  andMask = 64'b1111111111111111111111100000000000000000000000000000000000000000;
        6'd23:  andMask = 64'b1111111111111111111111110000000000000000000000000000000000000000;
        6'd24:  andMask = 64'b1111111111111111111111111000000000000000000000000000000000000000;
        6'd25:  andMask = 64'b1111111111111111111111111100000000000000000000000000000000000000;
        6'd26:  andMask = 64'b1111111111111111111111111110000000000000000000000000000000000000;
        6'd27:  andMask = 64'b1111111111111111111111111111000000000000000000000000000000000000;
        6'd28:  andMask = 64'b1111111111111111111111111111100000000000000000000000000000000000;
        6'd29:  andMask = 64'b1111111111111111111111111111110000000000000000000000000000000000;
        6'd30:  andMask = 64'b1111111111111111111111111111111000000000000000000000000000000000;
        6'd31:  andMask = 64'b1111111111111111111111111111111100000000000000000000000000000000;
        6'd32:  andMask = 64'b1111111111111111111111111111111110000000000000000000000000000000;
        6'd33:  andMask = 64'b1111111111111111111111111111111111000000000000000000000000000000;
        6'd34:  andMask = 64'b1111111111111111111111111111111111100000000000000000000000000000;
        6'd35:  andMask = 64'b1111111111111111111111111111111111110000000000000000000000000000;
        6'd36:  andMask = 64'b1111111111111111111111111111111111111000000000000000000000000000;
        6'd37:  andMask = 64'b1111111111111111111111111111111111111100000000000000000000000000;
        6'd38:  andMask = 64'b1111111111111111111111111111111111111110000000000000000000000000;
        6'd39:  andMask = 64'b1111111111111111111111111111111111111111000000000000000000000000;
        6'd40:  andMask = 64'b1111111111111111111111111111111111111111100000000000000000000000;
        6'd41:  andMask = 64'b1111111111111111111111111111111111111111110000000000000000000000;
        6'd42:  andMask = 64'b1111111111111111111111111111111111111111111000000000000000000000;
        6'd43:  andMask = 64'b1111111111111111111111111111111111111111111100000000000000000000;
        6'd44:  andMask = 64'b1111111111111111111111111111111111111111111110000000000000000000;
        6'd45:  andMask = 64'b1111111111111111111111111111111111111111111111000000000000000000;
        6'd46:  andMask = 64'b1111111111111111111111111111111111111111111111100000000000000000;
        6'd47:  andMask = 64'b1111111111111111111111111111111111111111111111110000000000000000;
        6'd48:  andMask = 64'b1111111111111111111111111111111111111111111111111000000000000000;
        6'd49:  andMask = 64'b1111111111111111111111111111111111111111111111111100000000000000;
        6'd50:  andMask = 64'b1111111111111111111111111111111111111111111111111110000000000000;
        6'd51:  andMask = 64'b1111111111111111111111111111111111111111111111111111000000000000;
        6'd52:  andMask = 64'b1111111111111111111111111111111111111111111111111111100000000000;
        6'd53:  andMask = 64'b1111111111111111111111111111111111111111111111111111110000000000;
        6'd54:  andMask = 64'b1111111111111111111111111111111111111111111111111111111000000000;
        6'd55:  andMask = 64'b1111111111111111111111111111111111111111111111111111111100000000;
        6'd56:  andMask = 64'b1111111111111111111111111111111111111111111111111111111110000000;
        6'd57:  andMask = 64'b1111111111111111111111111111111111111111111111111111111111000000;
        6'd58:  andMask = 64'b1111111111111111111111111111111111111111111111111111111111100000;
        6'd59:  andMask = 64'b1111111111111111111111111111111111111111111111111111111111110000;
        6'd60:  andMask = 64'b1111111111111111111111111111111111111111111111111111111111111000;
        6'd61:  andMask = 64'b1111111111111111111111111111111111111111111111111111111111111100;
        6'd62:  andMask = 64'b1111111111111111111111111111111111111111111111111111111111111110;
        6'd63:  andMask = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        default : andMask = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    endcase

    case( message_length[5:0])
        6'd0:   orMask = 64'b1000000000000000000000000000000000000000000000000000000000000000;
        6'd1:   orMask = 64'b0100000000000000000000000000000000000000000000000000000000000000;
        6'd2:   orMask = 64'b0010000000000000000000000000000000000000000000000000000000000000;
        6'd3:   orMask = 64'b0001000000000000000000000000000000000000000000000000000000000000;
        6'd4:   orMask = 64'b0000100000000000000000000000000000000000000000000000000000000000;
        6'd5:   orMask = 64'b0000010000000000000000000000000000000000000000000000000000000000;
        6'd6:   orMask = 64'b0000001000000000000000000000000000000000000000000000000000000000;
        6'd7:   orMask = 64'b0000000100000000000000000000000000000000000000000000000000000000;
        6'd8:   orMask = 64'b0000000010000000000000000000000000000000000000000000000000000000;
        6'd9:   orMask = 64'b0000000001000000000000000000000000000000000000000000000000000000;
        6'd10:  orMask = 64'b0000000000100000000000000000000000000000000000000000000000000000;
        6'd11:  orMask = 64'b0000000000010000000000000000000000000000000000000000000000000000;
        6'd12:  orMask = 64'b0000000000001000000000000000000000000000000000000000000000000000;
        6'd13:  orMask = 64'b0000000000000100000000000000000000000000000000000000000000000000;
        6'd14:  orMask = 64'b0000000000000010000000000000000000000000000000000000000000000000;
        6'd15:  orMask = 64'b0000000000000001000000000000000000000000000000000000000000000000;
        6'd16:  orMask = 64'b0000000000000000100000000000000000000000000000000000000000000000;
        6'd17:  orMask = 64'b0000000000000000010000000000000000000000000000000000000000000000;
        6'd18:  orMask = 64'b0000000000000000001000000000000000000000000000000000000000000000;
        6'd19:  orMask = 64'b0000000000000000000100000000000000000000000000000000000000000000;
        6'd20:  orMask = 64'b0000000000000000000010000000000000000000000000000000000000000000;
        6'd21:  orMask = 64'b0000000000000000000001000000000000000000000000000000000000000000;
        6'd22:  orMask = 64'b0000000000000000000000100000000000000000000000000000000000000000;
        6'd23:  orMask = 64'b0000000000000000000000010000000000000000000000000000000000000000;
        6'd24:  orMask = 64'b0000000000000000000000001000000000000000000000000000000000000000;
        6'd25:  orMask = 64'b0000000000000000000000000100000000000000000000000000000000000000;
        6'd26:  orMask = 64'b0000000000000000000000000010000000000000000000000000000000000000;
        6'd27:  orMask = 64'b0000000000000000000000000001000000000000000000000000000000000000;
        6'd28:  orMask = 64'b0000000000000000000000000000100000000000000000000000000000000000;
        6'd29:  orMask = 64'b0000000000000000000000000000010000000000000000000000000000000000;
        6'd30:  orMask = 64'b0000000000000000000000000000001000000000000000000000000000000000;
        6'd31:  orMask = 64'b0000000000000000000000000000000100000000000000000000000000000000;
        6'd32:  orMask = 64'b0000000000000000000000000000000010000000000000000000000000000000;
        6'd33:  orMask = 64'b0000000000000000000000000000000001000000000000000000000000000000;
        6'd34:  orMask = 64'b0000000000000000000000000000000000100000000000000000000000000000;
        6'd35:  orMask = 64'b0000000000000000000000000000000000010000000000000000000000000000;
        6'd36:  orMask = 64'b0000000000000000000000000000000000001000000000000000000000000000;
        6'd37:  orMask = 64'b0000000000000000000000000000000000000100000000000000000000000000;
        6'd38:  orMask = 64'b0000000000000000000000000000000000000010000000000000000000000000;
        6'd39:  orMask = 64'b0000000000000000000000000000000000000001000000000000000000000000;
        6'd40:  orMask = 64'b0000000000000000000000000000000000000000100000000000000000000000;
        6'd41:  orMask = 64'b0000000000000000000000000000000000000000010000000000000000000000;
        6'd42:  orMask = 64'b0000000000000000000000000000000000000000001000000000000000000000;
        6'd43:  orMask = 64'b0000000000000000000000000000000000000000000100000000000000000000;
        6'd44:  orMask = 64'b0000000000000000000000000000000000000000000010000000000000000000;
        6'd45:  orMask = 64'b0000000000000000000000000000000000000000000001000000000000000000;
        6'd46:  orMask = 64'b0000000000000000000000000000000000000000000000100000000000000000;
        6'd47:  orMask = 64'b0000000000000000000000000000000000000000000000010000000000000000;
        6'd48:  orMask = 64'b0000000000000000000000000000000000000000000000001000000000000000;
        6'd49:  orMask = 64'b0000000000000000000000000000000000000000000000000100000000000000;
        6'd50:  orMask = 64'b0000000000000000000000000000000000000000000000000010000000000000;
        6'd51:  orMask = 64'b0000000000000000000000000000000000000000000000000001000000000000;
        6'd52:  orMask = 64'b0000000000000000000000000000000000000000000000000000100000000000;
        6'd53:  orMask = 64'b0000000000000000000000000000000000000000000000000000010000000000;
        6'd54:  orMask = 64'b0000000000000000000000000000000000000000000000000000001000000000;
        6'd55:  orMask = 64'b0000000000000000000000000000000000000000000000000000000100000000;
        6'd56:  orMask = 64'b0000000000000000000000000000000000000000000000000000000010000000;
        6'd57:  orMask = 64'b0000000000000000000000000000000000000000000000000000000001000000;
        6'd58:  orMask = 64'b0000000000000000000000000000000000000000000000000000000000100000;
        6'd59:  orMask = 64'b0000000000000000000000000000000000000000000000000000000000010000;
        6'd60:  orMask = 64'b0000000000000000000000000000000000000000000000000000000000001000;
        6'd61:  orMask = 64'b0000000000000000000000000000000000000000000000000000000000000100;
        6'd62:  orMask = 64'b0000000000000000000000000000000000000000000000000000000000000010;
        6'd63:  orMask = 64'b0000000000000000000000000000000000000000000000000000000000000001;
        default : orMask = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    endcase
end
endmodule